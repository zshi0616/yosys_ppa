module sky130_fd_sc_lp__fa (
    COUT,  
    SUM,   
    A,     
    B,     
    CIN    
);
    output COUT; 
    output SUM;  
    input  A;    
    input  B;    
    input  CIN;  
    wire or0_out;      
    wire and0_out;     
    wire and1_out;     
    wire and2_out;     
    wire nor0_out;     
    wire nor1_out;     
    wire or1_out_COUT; 
    wire or2_out_SUM;  
    or  or0  (or0_out, CIN, B);
    and and0 (and0_out, or0_out, A);
    and and1 (and1_out, B, CIN);
    or  or1  (or1_out_COUT, and1_out, and0_out);
    buf buf0 (COUT, or1_out_COUT);
    and and2 (and2_out, CIN, A, B);
    nor nor0 (nor0_out, A, or0_out);
    nor nor1 (nor1_out, nor0_out, COUT);
    or  or2  (or2_out_SUM, nor1_out, and2_out);
    buf buf1 (SUM, or2_out_SUM);
endmodule
module design1 (MO, IN0, IN1, IN2, IN3, S);
   input IN0;
   input IN1;
   input IN2;
   input IN3;
   input [1:0] S;
   output MO;
   wire IN0_in;
   wire IN1_in;
   wire IN2_in;
   wire IN3_in;
   wire S1_in;
   wire S0_in;
   buf(IN0_in, IN0);
   buf(IN1_in, IN1);
   buf(IN2_in, IN2);
   buf(IN3_in, IN3);
   buf(S1_in, S[1]);
   buf(S0_in, S[0]);
   wire   tmp_MO;
   specify
      (IN0 => MO) = (0, 0);
      (IN1 => MO) = (0, 0);
      (IN2 => MO) = (0, 0);
      (IN3 => MO) = (0, 0);
      (S[1] => MO) = (0, 0);
      (S[0] => MO) = (0, 0);
   endspecify
   assign tmp_MO = S1_in ? (S0_in ? IN3_in : IN2_in) : (S0_in ? IN1_in : IN0_in);
   buf (MO, tmp_MO);
endmodule

module design2 (MO, IN0, IN1, IN2, IN3, S);
   input IN0;
   input IN1;
   input IN2;
   input IN3;
   input [1:0] S;
   output reg MO;

   always @(*)
     case(S)
       2'b00: MO = IN0;
       2'b01: MO = IN1;
       2'b10: MO = IN2;
       2'b11: MO = IN3;
     endcase
endmodule

module miter();
wire  MO1, MO2;
design1 inst1 (.MO(MO1),.IN0(IN0),.IN1(IN1),.IN2(IN2),.IN3(IN3),.S(S));
design2 inst2 (.MO(MO2),.IN0(IN0),.IN1(IN1),.IN2(IN2),.IN3(IN3),.S(S));
always @* begin
assert(MO1 == MO2);
end
endmodule